b0VIM 8.0      KaX@�#  kicodevs                                supertitan                              ~kicodevs/kuma-workspace/wasi-chrono/src/main.rs                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad  �	  �
     :       �  �  �  �  �  l  4  �  �  �  �  �  {  n  [  T  5    �  �  �  �  �  �  �  �  {  y  x  l  <    �  �  u  C          �  �  �  �  �  �  �  �  �  \  )  #  "    �
  �
  �
  �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   }}}     }         let ep = get_epoch(&Utc);     fn get_epoch_utc() {     #[test]      }         let ep = get_epoch(&FixedOffset::east(0));     fn get_epoch_fixed_offset_0() {     #[test]      }         let ep = get_epoch(&Local);     fn get_epoch_local() {     #[test]          use super::*; mod tests { #[cfg(test)]  }     println!("{:?}", as_uuid("te2".to_string()));     println!("{:?}", as_uuid("tet".to_string()));     println!("{:?}", get_epoch(&Local));     println!("{:?}", get_epoch(&FixedOffset::east(0)));     println!("{:?}", get_epoch(&FixedOffset::east(9 * 3600)));     println!("{:?}", get_epoch(&Utc));     println!("Hello, world! {}", Local::now()); fn main() {  }         timezone.ymd(1900, 1, 1).and_hms(0, 0, 0) {     T: TimeZone, where fn get_epoch<T>(timezone: &T) -> DateTime<T>  }     }         Err(_) => Uuid::nil(),         Ok(uuid) => uuid,     match Uuid::parse_str(s) {     };         s.as_str()     } else {         reconstructed.as_str()          }             reconstructed.push(c);         for c in s.chars().skip(1).take(s.len() - 2) {         // reconstruct the string without the braces     let s = if s.starts_with('{') && s.ends_with('}') {     let mut reconstructed = String::new(); pub(crate) fn as_uuid(s: String) -> Uuid {  use uuid::Uuid; //use chrono::Local; use chrono::prelude::*; 